//=================================================================================================
//  File Name    : Encoder.v
//  Description  : 
//      This module implements the C-PHY encoder, which generates the required 3-phase signal
//      levels (A, B, C) from a 3-bit symbol input. The encoder transitions between six valid
//      states (X+, X-, Y+, Y-, Z+, Z-) to represent encoded data through differential signaling.
//      These states are cycled through based on the symbol input using clockwise and counter-
//      clockwise rotation, with or without polarity inversion.
//
//      The output drive levels are generated by setting pull-up (PU) and pull-down (PD) control
//      signals for each phase. The module ensures proper electrical levels (VDD, GND, 0.5VDD)
//      through a tri-state buffer style control logic, avoiding short-circuit current during 
//      transitions.
//
//  Key Inputs    : 
//      - RstN            : Active-low reset
//      - EncoderEn       : Enable signal for the encoder operation
//      - TxSymbolClkHS   : High-speed clock for symbol processing
//      - Sym             : 3-bit input symbol to be encoded
//
//  Key Outputs   : 
//      - A, B, C         : 2-bit (PU, PD) encoded output signals representing the three C-PHY phases
//
//  Author       : Youssef Ehab
//  Date         : 10/5/2025
//=================================================================================================

module Encoder(
    input            RstN,
    input            EncoderEn,
    input            TxSymbolClkHS,
    input      [2:0] Sym,
    output wire [1:0] A,
    output wire [1:0] B,
    output wire [1:0] C
);

reg [2:0] State;
reg [2:0] State_Intermediate;
reg       PU_A_Intermediate;
reg       PD_A_Intermediate;
reg       PU_B_Intermediate;
reg       PD_B_Intermediate;
reg       PU_C_Intermediate;
reg       PD_C_Intermediate;

reg  PU_A,PD_A,PU_B,PD_B,PU_C,PD_C;


// Concatenate into 2-bit signals
           assign A = {PU_A, PD_A};
           assign B = {PU_B, PD_B};
           assign C = {PU_C, PD_C};

always @(posedge TxSymbolClkHS, negedge RstN) begin
    if(!RstN) begin
        State <= 3'b100;
        PU_A <= 1'b0;
        PD_A <= 1'b1;
        PU_B <= 1'b0;
        PD_B <= 1'b1;
        PU_C <= 1'b0;
        PD_C <= 1'b1;
        //Reset value is set to one to drive zero volatge on the tri-State buffers to avoid short circuit currents
    end
    else begin
        if(EncoderEn) begin

            PU_A <= PU_A_Intermediate;
            PD_A <= PD_A_Intermediate;
            PU_B <= PU_B_Intermediate;
            PD_B <= PD_B_Intermediate;
            PU_C <= PU_C_Intermediate;
            PD_C <= PD_C_Intermediate;

            State <= State_Intermediate;

        end
        else begin
            State <= 3'b100;
            PU_A <= 1'b0;
            PD_A <= 1'b1;
            PU_B <= 1'b0;
            PD_B <= 1'b1;
            PU_C <= 1'b0;
            PD_C <= 1'b1;
            //Reset value is set to one to drive zero volatge on the tri-State buffers to avoid short circuit currents
        end
    end
end


//for the circuit to give vdd     : PU = 1 , PD = 0
//for the circuit to give 0       : PU = 0 , PD = 1
//for the circuit to give 0.5*vdd : PU = 1 , PD = 1

always @(*) begin

    case(State)
        3'b100: begin     //X+
            PU_A_Intermediate = 1'b1;
            PD_A_Intermediate = 1'b0;
            PU_B_Intermediate = 1'b0;
            PD_B_Intermediate = 1'b1;
            PU_C_Intermediate = 1'b1;
            PD_C_Intermediate = 1'b1;
        end
        3'b011: begin     //X-
            PU_A_Intermediate = 1'b0;
            PD_A_Intermediate = 1'b1;
            PU_B_Intermediate = 1'b1;
            PD_B_Intermediate = 1'b0;
            PU_C_Intermediate = 1'b1;
            PD_C_Intermediate = 1'b1;
        end
        3'b010: begin     //Y+
            PU_A_Intermediate = 1'b1;
            PD_A_Intermediate = 1'b1;
            PU_B_Intermediate = 1'b1;
            PD_B_Intermediate = 1'b0;
            PU_C_Intermediate = 1'b0;
            PD_C_Intermediate = 1'b1;
        end
        3'b101: begin     //Y-
            PU_A_Intermediate = 1'b1;
            PD_A_Intermediate = 1'b1;
            PU_B_Intermediate = 1'b0;
            PD_B_Intermediate = 1'b1;
            PU_C_Intermediate = 1'b1;
            PD_C_Intermediate = 1'b0;
        end
        3'b001: begin     //Z+
            PU_A_Intermediate = 1'b0;
            PD_A_Intermediate = 1'b1;
            PU_B_Intermediate = 1'b1;
            PD_B_Intermediate = 1'b1;
            PU_C_Intermediate = 1'b1;
            PD_C_Intermediate = 1'b0;
        end
        3'b110: begin     //Z-
            PU_A_Intermediate = 1'b1;
            PD_A_Intermediate = 1'b0;
            PU_B_Intermediate = 1'b1;
            PD_B_Intermediate = 1'b1;
            PU_C_Intermediate = 1'b0;
            PD_C_Intermediate = 1'b1;
        end
        default: begin     
            PU_A_Intermediate = 1'b0;
            PD_A_Intermediate = 1'b1;
            PU_B_Intermediate = 1'b0;
            PD_B_Intermediate = 1'b1;
            PU_C_Intermediate = 1'b0;
            PD_C_Intermediate = 1'b1;
        end
    endcase

    case(Sym)
        3'b000:  State_Intermediate = {State[1:0],State[2]};  //Rotate CCW, Same Polarity
        3'b001:  State_Intermediate = ~{State[1:0],State[2]}; //Rotate CCW, Opposite Polarity
        3'b010:  State_Intermediate = {State[0],State[2:1]};  //Rotate CW,  Same Polarity
        3'b011:  State_Intermediate = ~{State[0],State[2:1]}; //Rotate CW,  Opposite Polarity
        3'b100:  State_Intermediate = ~State;                 //Same phase, Opposite polarity
        3'b101:  State_Intermediate = ~State;                 //Same phase, Opposite polarity
        3'b110:  State_Intermediate = ~State;                 //Same phase, Opposite polarity
        3'b111:  State_Intermediate = ~State;                 //Same phase, Opposite polarity
        default: State_Intermediate = State;
    endcase
end

endmodule